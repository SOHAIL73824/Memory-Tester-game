module tb_timer();
reg clock,rst;
reg decrement,load,stop;
reg [3:0] reconfig2;
reg [7:0] input_num;
wire time_stop;
wire [3:0] timedig1,timedig2;
wire outpulse,borrow,stop_upstream;


two_digit_timer testtime(clock,rst,stop,decrement,load,reconfig2,input_num,time_stop,timedig1,timedig2,outpulse,borrow,stop_upstream);
always
begin
 clock=0;
 #10;
 clock=1;
 #10;
end

initial 
begin
rst=0;
@(posedge clock);
#5 rst=1;stop=1;
@(posedge clock);
input_num=8'b00110011;
@(posedge clock);
#5 load=1;
@(posedge clock);
#5 load=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 decrement=1;
@(posedge clock);
#5 decrement=0;




end
endmodule
