`timescale 1ps/1ps
module tb_score();
reg clock,rst,green_user,auth_bit,win,loose,disp_button,log_out;
reg [3:0] level_num;
reg [2:0] internal_id;
wire [7:0] disp_out;
wire green_max;
integer i;

score_table test_score(clock,rst,log_out,green_user,internal_id,auth_bit,win,loose,disp_button,level_num,disp_out,green_max);
always
begin
 clock=0;
 #10;
 clock=1;
 #10;
end
 
initial 
begin
rst=0;
@(posedge clock);
#5 rst=1;log_out=0;
@(posedge clock);
#5 green_user=1; internal_id=3'b101;disp_button=1;
@(posedge clock);
#5 auth_bit=1;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0001;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0010;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0011;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0100;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0101;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0001;
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 loose=1;
@(posedge clock);
#5 loose=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 log_out=1;
@(posedge clock);
#5 log_out=0;

//green_max
@(posedge clock);
#5 green_user=1; internal_id=3'b110;disp_button=1;
@(posedge clock);
#5 auth_bit=1;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0001;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0010;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0011;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0100;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0101;
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0001;
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 level_num=4'b0010;
@(posedge clock);
#5 win=1;
@(posedge clock);
#5 win=0;
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
@(posedge clock);
#5 log_out=1;
@(posedge clock);
#5 log_out=0;

end

endmodule
